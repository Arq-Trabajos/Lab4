module ej (
    input [1:0] ALUControl, input [31:0] A, input [31:0] B, input [31:0] Sum,
    output [3:0] ALUFlags, output [31:0] result
);

endmodule

module mux4_1(
    input [1:0] S, input A, B, C, D,
    output O
);
    
endmodule